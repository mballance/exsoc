/****************************************************************************
 * axi_slave.sv
 ****************************************************************************/

/**
 * Module: axi_slave
 * 
 * TODO: Add module documentation
 */
module axi_slave(
		input			clk,
		input			reset,
		axi4_if.aw_slave		aw_1,
		axi4_if.b_slave			b_1,
		axi4_if.ar_slave		ar_1,
		axi4_if.r_slave			r_1);


endmodule

