
module top;

	reg clk, rst;

	axi4_if axi(clk, rst);

endmodule

